LEDCUBE
C2 1 3 1µF IC=0
C1 37 0 1µF IC=0
R4 7 6 1k
C3 1 2 1µF IC=0
R2 31 10 1k
R3 9 8 1k
R5 5 4 1k
R1 37 1 220

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
